module andgate (A, B, F);

//inputs
input A;
input B;

//outputs
output F;

assign F = A & B;

endmodule